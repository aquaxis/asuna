/*
 * Copyright (C)2005-2024 AQUAXIS TECHNOLOGY.
 *  Don't remove this header.
 * When you use this source, there is a need to inherit this header.
 *
 * This software is released under the MIT License.
 * https://opensource.org/license/mit
 */

 module aq_div31x31(
	input			RST_N,
	input			CLK,
	input [30:0]	DINA,
	input [30:0]	DINB,
	output [30:0]	QOUT,
	output [30:0]	ROUT
);
reg [62:0] r00r;
reg [62:0] r01r;
reg [62:0] r02r;
reg [62:0] r03r;
reg [62:0] r04r;
reg [62:0] r05r;
reg [62:0] r06r;
reg [62:0] r07r;
reg [62:0] r08r;
reg [62:0] r09r;
reg [62:0] r10r;
reg [62:0] r11r;
reg [62:0] r12r;
reg [62:0] r13r;
reg [62:0] r14r;
reg [62:0] r15r;
reg [62:0] r16r;
reg [62:0] r17r;
reg [62:0] r18r;
reg [62:0] r19r;
reg [62:0] r20r;
reg [62:0] r21r;
reg [62:0] r22r;
reg [62:0] r23r;
reg [62:0] r24r;
reg [62:0] r25r;
reg [62:0] r26r;
reg [62:0] r27r;
reg [62:0] r28r;
reg [62:0] r29r;
reg [62:0] r30r;
reg [62:0] r31r;
reg [30:0] s00r;
reg [30:0] s01r;
reg [30:0] s02r;
reg [30:0] s03r;
reg [30:0] s04r;
reg [30:0] s05r;
reg [30:0] s06r;
reg [30:0] s07r;
reg [30:0] s08r;
reg [30:0] s09r;
reg [30:0] s10r;
reg [30:0] s11r;
reg [30:0] s12r;
reg [30:0] s13r;
reg [30:0] s14r;
reg [30:0] s15r;
reg [30:0] s16r;
reg [30:0] s17r;
reg [30:0] s18r;
reg [30:0] s19r;
reg [30:0] s20r;
reg [30:0] s21r;
reg [30:0] s22r;
reg [30:0] s23r;
reg [30:0] s24r;
reg [30:0] s25r;
reg [30:0] s26r;
reg [30:0] s27r;
reg [30:0] s28r;
reg [30:0] s29r;
reg [30:0] s30r;
reg [30:0] s31r;
always @(negedge RST_N or posedge CLK) begin
	if(!RST_N) begin
		r00r <= 63'd0;
		r01r <= 63'd0;
		r02r <= 63'd0;
		r03r <= 63'd0;
		r04r <= 63'd0;
		r05r <= 63'd0;
		r06r <= 63'd0;
		r07r <= 63'd0;
		r08r <= 63'd0;
		r09r <= 63'd0;
		r10r <= 63'd0;
		r11r <= 63'd0;
		r12r <= 63'd0;
		r13r <= 63'd0;
		r14r <= 63'd0;
		r15r <= 63'd0;
		r16r <= 63'd0;
		r17r <= 63'd0;
		r18r <= 63'd0;
		r19r <= 63'd0;
		r20r <= 63'd0;
		r21r <= 63'd0;
		r22r <= 63'd0;
		r23r <= 63'd0;
		r24r <= 63'd0;
		r25r <= 63'd0;
		r26r <= 63'd0;
		r27r <= 63'd0;
		r28r <= 63'd0;
		r29r <= 63'd0;
		r30r <= 63'd0;
		r31r <= 63'd0;
		s00r <= 31'd0;
		s01r <= 31'd0;
		s02r <= 31'd0;
		s03r <= 31'd0;
		s04r <= 31'd0;
		s05r <= 31'd0;
		s06r <= 31'd0;
		s07r <= 31'd0;
		s08r <= 31'd0;
		s09r <= 31'd0;
		s10r <= 31'd0;
		s11r <= 31'd0;
		s12r <= 31'd0;
		s13r <= 31'd0;
		s14r <= 31'd0;
		s15r <= 31'd0;
		s16r <= 31'd0;
		s17r <= 31'd0;
		s18r <= 31'd0;
		s19r <= 31'd0;
		s20r <= 31'd0;
		s21r <= 31'd0;
		s22r <= 31'd0;
		s23r <= 31'd0;
		s24r <= 31'd0;
		s25r <= 31'd0;
		s26r <= 31'd0;
		s27r <= 31'd0;
		s28r <= 31'd0;
		s29r <= 31'd0;
		s30r <= 31'd0;
	end else begin
		// Stage: buffer
		r00r[62:0]	<= {1'b1, 31'd0, DINA};
		s00r 		<= DINB;

		// State: 01
		r01r[62:30]	<= ({1'b1,r00r[61:30]}) + (~{2'b00,s00r}) + 1;
		r01r[29:0]	<= r00r[29:0] ;
		s01r <= s00r;

		// State: 02
		r02r[61:29]	<= ({r01r[62],r01r[60:29]}) + (({33{r01r[62]}}^{2'b00,s01r}) + r01r[62]);
		r02r[62:62]	<= r01r[62:62] ;
		r02r[28:0]	<= r01r[28:0] ;
		s02r <= s01r;

		// State: 03
		r03r[60:28]	<= ({r02r[61],r02r[59:28]}) + (({33{r02r[61]}}^{2'b00,s02r}) + r02r[61]);
		r03r[62:61]	<= r02r[62:61] ;
		r03r[27:0]	<= r02r[27:0] ;
		s03r <= s02r;

		// State: 04
		r04r[59:27]	<= ({r03r[60],r03r[58:27]}) + (({33{r03r[60]}}^{2'b00,s03r}) + r03r[60]);
		r04r[62:60]	<= r03r[62:60] ;
		r04r[26:0]	<= r03r[26:0] ;
		s04r <= s03r;

		// State: 05
		r05r[58:26]	<= ({r04r[59],r04r[57:26]}) + (({33{r04r[59]}}^{2'b00,s04r}) + r04r[59]);
		r05r[62:59]	<= r04r[62:59] ;
		r05r[25:0]	<= r04r[25:0] ;
		s05r <= s04r;

		// State: 06
		r06r[57:25]	<= ({r05r[58],r05r[56:25]}) + (({33{r05r[58]}}^{2'b00,s05r}) + r05r[58]);
		r06r[62:58]	<= r05r[62:58] ;
		r06r[24:0]	<= r05r[24:0] ;
		s06r <= s05r;

		// State: 07
		r07r[56:24]	<= ({r06r[57],r06r[55:24]}) + (({33{r06r[57]}}^{2'b00,s06r}) + r06r[57]);
		r07r[62:57]	<= r06r[62:57] ;
		r07r[23:0]	<= r06r[23:0] ;
		s07r <= s06r;

		// State: 08
		r08r[55:23]	<= ({r07r[56],r07r[54:23]}) + (({33{r07r[56]}}^{2'b00,s07r}) + r07r[56]);
		r08r[62:56]	<= r07r[62:56] ;
		r08r[22:0]	<= r07r[22:0] ;
		s08r <= s07r;

		// State: 09
		r09r[54:22]	<= ({r08r[55],r08r[53:22]}) + (({33{r08r[55]}}^{2'b00,s08r}) + r08r[55]);
		r09r[62:55]	<= r08r[62:55] ;
		r09r[21:0]	<= r08r[21:0] ;
		s09r <= s08r;

		// State: 10
		r10r[53:21]	<= ({r09r[54],r09r[52:21]}) + (({33{r09r[54]}}^{2'b00,s09r}) + r09r[54]);
		r10r[62:54]	<= r09r[62:54] ;
		r10r[20:0]	<= r09r[20:0] ;
		s10r <= s09r;

		// State: 11
		r11r[52:20]	<= ({r10r[53],r10r[51:20]}) + (({33{r10r[53]}}^{2'b00,s10r}) + r10r[53]);
		r11r[62:53]	<= r10r[62:53] ;
		r11r[19:0]	<= r10r[19:0] ;
		s11r <= s10r;

		// State: 12
		r12r[51:19]	<= ({r11r[52],r11r[50:19]}) + (({33{r11r[52]}}^{2'b00,s11r}) + r11r[52]);
		r12r[62:52]	<= r11r[62:52] ;
		r12r[18:0]	<= r11r[18:0] ;
		s12r <= s11r;

		// State: 13
		r13r[50:18]	<= ({r12r[51],r12r[49:18]}) + (({33{r12r[51]}}^{2'b00,s12r}) + r12r[51]);
		r13r[62:51]	<= r12r[62:51] ;
		r13r[17:0]	<= r12r[17:0] ;
		s13r <= s12r;

		// State: 14
		r14r[49:17]	<= ({r13r[50],r13r[48:17]}) + (({33{r13r[50]}}^{2'b00,s13r}) + r13r[50]);
		r14r[62:50]	<= r13r[62:50] ;
		r14r[16:0]	<= r13r[16:0] ;
		s14r <= s13r;

		// State: 15
		r15r[48:16]	<= ({r14r[49],r14r[47:16]}) + (({33{r14r[49]}}^{2'b00,s14r}) + r14r[49]);
		r15r[62:49]	<= r14r[62:49] ;
		r15r[15:0]	<= r14r[15:0] ;
		s15r <= s14r;

		// State: 16
		r16r[47:15]	<= ({r15r[48],r15r[46:15]}) + (({33{r15r[48]}}^{2'b00,s15r}) + r15r[48]);
		r16r[62:48]	<= r15r[62:48] ;
		r16r[14:0]	<= r15r[14:0] ;
		s16r <= s15r;

		// State: 17
		r17r[46:14]	<= ({r16r[47],r16r[45:14]}) + (({33{r16r[47]}}^{2'b00,s16r}) + r16r[47]);
		r17r[62:47]	<= r16r[62:47] ;
		r17r[13:0]	<= r16r[13:0] ;
		s17r <= s16r;

		// State: 18
		r18r[45:13]	<= ({r17r[46],r17r[44:13]}) + (({33{r17r[46]}}^{2'b00,s17r}) + r17r[46]);
		r18r[62:46]	<= r17r[62:46] ;
		r18r[12:0]	<= r17r[12:0] ;
		s18r <= s17r;

		// State: 19
		r19r[44:12]	<= ({r18r[45],r18r[43:12]}) + (({33{r18r[45]}}^{2'b00,s18r}) + r18r[45]);
		r19r[62:45]	<= r18r[62:45] ;
		r19r[11:0]	<= r18r[11:0] ;
		s19r <= s18r;

		// State: 20
		r20r[43:11]	<= ({r19r[44],r19r[42:11]}) + (({33{r19r[44]}}^{2'b00,s19r}) + r19r[44]);
		r20r[62:44]	<= r19r[62:44] ;
		r20r[10:0]	<= r19r[10:0] ;
		s20r <= s19r;

		// State: 21
		r21r[42:10]	<= ({r20r[43],r20r[41:10]}) + (({33{r20r[43]}}^{2'b00,s20r}) + r20r[43]);
		r21r[62:43]	<= r20r[62:43] ;
		r21r[9:0]	<= r20r[9:0] ;
		s21r <= s20r;

		// State: 22
		r22r[41:9]	<= ({r21r[42],r21r[40:9]}) + (({33{r21r[42]}}^{2'b00,s21r}) + r21r[42]);
		r22r[62:42]	<= r21r[62:42] ;
		r22r[8:0]	<= r21r[8:0] ;
		s22r <= s21r;

		// State: 23
		r23r[40:8]	<= ({r22r[41],r22r[39:8]}) + (({33{r22r[41]}}^{2'b00,s22r}) + r22r[41]);
		r23r[62:41]	<= r22r[62:41] ;
		r23r[7:0]	<= r22r[7:0] ;
		s23r <= s22r;

		// State: 24
		r24r[39:7]	<= ({r23r[40],r23r[38:7]}) + (({33{r23r[40]}}^{2'b00,s23r}) + r23r[40]);
		r24r[62:40]	<= r23r[62:40] ;
		r24r[6:0]	<= r23r[6:0] ;
		s24r <= s23r;

		// State: 25
		r25r[38:6]	<= ({r24r[39],r24r[37:6]}) + (({33{r24r[39]}}^{2'b00,s24r}) + r24r[39]);
		r25r[62:39]	<= r24r[62:39] ;
		r25r[5:0]	<= r24r[5:0] ;
		s25r <= s24r;

		// State: 26
		r26r[37:5]	<= ({r25r[38],r25r[36:5]}) + (({33{r25r[38]}}^{2'b00,s25r}) + r25r[38]);
		r26r[62:38]	<= r25r[62:38] ;
		r26r[4:0]	<= r25r[4:0] ;
		s26r <= s25r;

		// State: 27
		r27r[36:4]	<= ({r26r[37],r26r[35:4]}) + (({33{r26r[37]}}^{2'b00,s26r}) + r26r[37]);
		r27r[62:37]	<= r26r[62:37] ;
		r27r[3:0]	<= r26r[3:0] ;
		s27r <= s26r;

		// State: 28
		r28r[35:3]	<= ({r27r[36],r27r[34:3]}) + (({33{r27r[36]}}^{2'b00,s27r}) + r27r[36]);
		r28r[62:36]	<= r27r[62:36] ;
		r28r[2:0]	<= r27r[2:0] ;
		s28r <= s27r;

		// State: 29
		r29r[34:2]	<= ({r28r[35],r28r[33:2]}) + (({33{r28r[35]}}^{2'b00,s28r}) + r28r[35]);
		r29r[62:35]	<= r28r[62:35] ;
		r29r[1:0]	<= r28r[1:0] ;
		s29r <= s28r;

		// State: 30
		r30r[33:1]	<= ({r29r[34],r29r[32:1]}) + (({33{r29r[34]}}^{2'b00,s29r}) + r29r[34]);
		r30r[62:34]	<= r29r[62:34] ;
		r30r[0:0]	<= r29r[0:0] ;
		s30r <= s29r;

		// State: 31
		r31r[32:0]	<= ({r30r[33],r30r[31:0]}) + (({33{r30r[33]}}^{2'b00,s30r}) + r30r[33]);
		r31r[62:33]	<= r30r[62:33] ;
		s31r <= s30r;

	end
end
assign QOUT = r31r[62:32];
assign ROUT = (r31r[31])?(r31r[30:0]+s31r):r31r[30:0];
endmodule
