/*
 * Copyright (C)2005-2024 AQUAXIS TECHNOLOGY.
 *  Don't remove this header.
 * When you use this source, there is a need to inherit this header.
 *
 * This software is released under the MIT License.
 * https://opensource.org/license/mit
 */
 module aq_div32x32(
	input			RST_N,
	input			CLK,
	input [31:0]	DINA,
	input [31:0]	DINB,
	output [31:0]	DOUT
);
reg [64:0] r00r;
reg [64:0] r01r;
reg [64:0] r02r;
reg [64:0] r03r;
reg [64:0] r04r;
reg [64:0] r05r;
reg [64:0] r06r;
reg [64:0] r07r;
reg [64:0] r08r;
reg [64:0] r09r;
reg [64:0] r10r;
reg [64:0] r11r;
reg [64:0] r12r;
reg [64:0] r13r;
reg [64:0] r14r;
reg [64:0] r15r;
reg [64:0] r16r;
reg [64:0] r17r;
reg [64:0] r18r;
reg [64:0] r19r;
reg [64:0] r20r;
reg [64:0] r21r;
reg [64:0] r22r;
reg [64:0] r23r;
reg [64:0] r24r;
reg [64:0] r25r;
reg [64:0] r26r;
reg [64:0] r27r;
reg [64:0] r28r;
reg [64:0] r29r;
reg [64:0] r30r;
reg [64:0] r31r;
reg [64:0] r32r;
reg [31:0] s00r;
reg [31:0] s01r;
reg [31:0] s02r;
reg [31:0] s03r;
reg [31:0] s04r;
reg [31:0] s05r;
reg [31:0] s06r;
reg [31:0] s07r;
reg [31:0] s08r;
reg [31:0] s09r;
reg [31:0] s10r;
reg [31:0] s11r;
reg [31:0] s12r;
reg [31:0] s13r;
reg [31:0] s14r;
reg [31:0] s15r;
reg [31:0] s16r;
reg [31:0] s17r;
reg [31:0] s18r;
reg [31:0] s19r;
reg [31:0] s20r;
reg [31:0] s21r;
reg [31:0] s22r;
reg [31:0] s23r;
reg [31:0] s24r;
reg [31:0] s25r;
reg [31:0] s26r;
reg [31:0] s27r;
reg [31:0] s28r;
reg [31:0] s29r;
reg [31:0] s30r;
reg [31:0] s31r;
always @(negedge RST_N or posedge CLK) begin
	if(!RST_N) begin
		r00r <= 65'd0;
		r01r <= 65'd0;
		r02r <= 65'd0;
		r03r <= 65'd0;
		r04r <= 65'd0;
		r05r <= 65'd0;
		r06r <= 65'd0;
		r07r <= 65'd0;
		r08r <= 65'd0;
		r09r <= 65'd0;
		r10r <= 65'd0;
		r11r <= 65'd0;
		r12r <= 65'd0;
		r13r <= 65'd0;
		r14r <= 65'd0;
		r15r <= 65'd0;
		r16r <= 65'd0;
		r17r <= 65'd0;
		r18r <= 65'd0;
		r19r <= 65'd0;
		r20r <= 65'd0;
		r21r <= 65'd0;
		r22r <= 65'd0;
		r23r <= 65'd0;
		r24r <= 65'd0;
		r25r <= 65'd0;
		r26r <= 65'd0;
		r27r <= 65'd0;
		r28r <= 65'd0;
		r29r <= 65'd0;
		r30r <= 65'd0;
		r31r <= 65'd0;
		r32r <= 65'd0;
		s00r <= 32'd0;
		s01r <= 32'd0;
		s02r <= 32'd0;
		s03r <= 32'd0;
		s04r <= 32'd0;
		s05r <= 32'd0;
		s06r <= 32'd0;
		s07r <= 32'd0;
		s08r <= 32'd0;
		s09r <= 32'd0;
		s10r <= 32'd0;
		s11r <= 32'd0;
		s12r <= 32'd0;
		s13r <= 32'd0;
		s14r <= 32'd0;
		s15r <= 32'd0;
		s16r <= 32'd0;
		s17r <= 32'd0;
		s18r <= 32'd0;
		s19r <= 32'd0;
		s20r <= 32'd0;
		s21r <= 32'd0;
		s22r <= 32'd0;
		s23r <= 32'd0;
		s24r <= 32'd0;
		s25r <= 32'd0;
		s26r <= 32'd0;
		s27r <= 32'd0;
		s28r <= 32'd0;
		s29r <= 32'd0;
		s30r <= 32'd0;
		s31r <= 32'd0;
	end else begin
		// Stage: buffer
		r00r[64:0]	<= {1'b1, 32'd0, DINA};
		s00r 		<= DINB;

		// State: 01
		r01r[64:31]	<= ({1'b1,r00r[63:31]}) + (~{2'b00,s00r}) + 1;
		r01r[30:0]	<= r00r[30:0] ;
		s01r <= s00r;

		// State: 02
		r02r[63:30]	<= ({r01r[64],r01r[62:30]}) + (({34{r01r[64]}}^{2'b00,s01r}) + r01r[64]);
		r02r[64:64]	<= r01r[64:64] ;
		r02r[29:0]	<= r01r[29:0] ;
		s02r <= s01r;

		// State: 03
		r03r[62:29]	<= ({r02r[63],r02r[61:29]}) + (({34{r02r[63]}}^{2'b00,s02r}) + r02r[63]);
		r03r[64:63]	<= r02r[64:63] ;
		r03r[28:0]	<= r02r[28:0] ;
		s03r <= s02r;

		// State: 04
		r04r[61:28]	<= ({r03r[62],r03r[60:28]}) + (({34{r03r[62]}}^{2'b00,s03r}) + r03r[62]);
		r04r[64:62]	<= r03r[64:62] ;
		r04r[27:0]	<= r03r[27:0] ;
		s04r <= s03r;

		// State: 05
		r05r[60:27]	<= ({r04r[61],r04r[59:27]}) + (({34{r04r[61]}}^{2'b00,s04r}) + r04r[61]);
		r05r[64:61]	<= r04r[64:61] ;
		r05r[26:0]	<= r04r[26:0] ;
		s05r <= s04r;

		// State: 06
		r06r[59:26]	<= ({r05r[60],r05r[58:26]}) + (({34{r05r[60]}}^{2'b00,s05r}) + r05r[60]);
		r06r[64:60]	<= r05r[64:60] ;
		r06r[25:0]	<= r05r[25:0] ;
		s06r <= s05r;

		// State: 07
		r07r[58:25]	<= ({r06r[59],r06r[57:25]}) + (({34{r06r[59]}}^{2'b00,s06r}) + r06r[59]);
		r07r[64:59]	<= r06r[64:59] ;
		r07r[24:0]	<= r06r[24:0] ;
		s07r <= s06r;

		// State: 08
		r08r[57:24]	<= ({r07r[58],r07r[56:24]}) + (({34{r07r[58]}}^{2'b00,s07r}) + r07r[58]);
		r08r[64:58]	<= r07r[64:58] ;
		r08r[23:0]	<= r07r[23:0] ;
		s08r <= s07r;

		// State: 09
		r09r[56:23]	<= ({r08r[57],r08r[55:23]}) + (({34{r08r[57]}}^{2'b00,s08r}) + r08r[57]);
		r09r[64:57]	<= r08r[64:57] ;
		r09r[22:0]	<= r08r[22:0] ;
		s09r <= s08r;

		// State: 10
		r10r[55:22]	<= ({r09r[56],r09r[54:22]}) + (({34{r09r[56]}}^{2'b00,s09r}) + r09r[56]);
		r10r[64:56]	<= r09r[64:56] ;
		r10r[21:0]	<= r09r[21:0] ;
		s10r <= s09r;

		// State: 11
		r11r[54:21]	<= ({r10r[55],r10r[53:21]}) + (({34{r10r[55]}}^{2'b00,s10r}) + r10r[55]);
		r11r[64:55]	<= r10r[64:55] ;
		r11r[20:0]	<= r10r[20:0] ;
		s11r <= s10r;

		// State: 12
		r12r[53:20]	<= ({r11r[54],r11r[52:20]}) + (({34{r11r[54]}}^{2'b00,s11r}) + r11r[54]);
		r12r[64:54]	<= r11r[64:54] ;
		r12r[19:0]	<= r11r[19:0] ;
		s12r <= s11r;

		// State: 13
		r13r[52:19]	<= ({r12r[53],r12r[51:19]}) + (({34{r12r[53]}}^{2'b00,s12r}) + r12r[53]);
		r13r[64:53]	<= r12r[64:53] ;
		r13r[18:0]	<= r12r[18:0] ;
		s13r <= s12r;

		// State: 14
		r14r[51:18]	<= ({r13r[52],r13r[50:18]}) + (({34{r13r[52]}}^{2'b00,s13r}) + r13r[52]);
		r14r[64:52]	<= r13r[64:52] ;
		r14r[17:0]	<= r13r[17:0] ;
		s14r <= s13r;

		// State: 15
		r15r[50:17]	<= ({r14r[51],r14r[49:17]}) + (({34{r14r[51]}}^{2'b00,s14r}) + r14r[51]);
		r15r[64:51]	<= r14r[64:51] ;
		r15r[16:0]	<= r14r[16:0] ;
		s15r <= s14r;

		// State: 16
		r16r[49:16]	<= ({r15r[50],r15r[48:16]}) + (({34{r15r[50]}}^{2'b00,s15r}) + r15r[50]);
		r16r[64:50]	<= r15r[64:50] ;
		r16r[15:0]	<= r15r[15:0] ;
		s16r <= s15r;

		// State: 17
		r17r[48:15]	<= ({r16r[49],r16r[47:15]}) + (({34{r16r[49]}}^{2'b00,s16r}) + r16r[49]);
		r17r[64:49]	<= r16r[64:49] ;
		r17r[14:0]	<= r16r[14:0] ;
		s17r <= s16r;

		// State: 18
		r18r[47:14]	<= ({r17r[48],r17r[46:14]}) + (({34{r17r[48]}}^{2'b00,s17r}) + r17r[48]);
		r18r[64:48]	<= r17r[64:48] ;
		r18r[13:0]	<= r17r[13:0] ;
		s18r <= s17r;

		// State: 19
		r19r[46:13]	<= ({r18r[47],r18r[45:13]}) + (({34{r18r[47]}}^{2'b00,s18r}) + r18r[47]);
		r19r[64:47]	<= r18r[64:47] ;
		r19r[12:0]	<= r18r[12:0] ;
		s19r <= s18r;

		// State: 20
		r20r[45:12]	<= ({r19r[46],r19r[44:12]}) + (({34{r19r[46]}}^{2'b00,s19r}) + r19r[46]);
		r20r[64:46]	<= r19r[64:46] ;
		r20r[11:0]	<= r19r[11:0] ;
		s20r <= s19r;

		// State: 21
		r21r[44:11]	<= ({r20r[45],r20r[43:11]}) + (({34{r20r[45]}}^{2'b00,s20r}) + r20r[45]);
		r21r[64:45]	<= r20r[64:45] ;
		r21r[10:0]	<= r20r[10:0] ;
		s21r <= s20r;

		// State: 22
		r22r[43:10]	<= ({r21r[44],r21r[42:10]}) + (({34{r21r[44]}}^{2'b00,s21r}) + r21r[44]);
		r22r[64:44]	<= r21r[64:44] ;
		r22r[9:0]	<= r21r[9:0] ;
		s22r <= s21r;

		// State: 23
		r23r[42:9]	<= ({r22r[43],r22r[41:9]}) + (({34{r22r[43]}}^{2'b00,s22r}) + r22r[43]);
		r23r[64:43]	<= r22r[64:43] ;
		r23r[8:0]	<= r22r[8:0] ;
		s23r <= s22r;

		// State: 24
		r24r[41:8]	<= ({r23r[42],r23r[40:8]}) + (({34{r23r[42]}}^{2'b00,s23r}) + r23r[42]);
		r24r[64:42]	<= r23r[64:42] ;
		r24r[7:0]	<= r23r[7:0] ;
		s24r <= s23r;

		// State: 25
		r25r[40:7]	<= ({r24r[41],r24r[39:7]}) + (({34{r24r[41]}}^{2'b00,s24r}) + r24r[41]);
		r25r[64:41]	<= r24r[64:41] ;
		r25r[6:0]	<= r24r[6:0] ;
		s25r <= s24r;

		// State: 26
		r26r[39:6]	<= ({r25r[40],r25r[38:6]}) + (({34{r25r[40]}}^{2'b00,s25r}) + r25r[40]);
		r26r[64:40]	<= r25r[64:40] ;
		r26r[5:0]	<= r25r[5:0] ;
		s26r <= s25r;

		// State: 27
		r27r[38:5]	<= ({r26r[39],r26r[37:5]}) + (({34{r26r[39]}}^{2'b00,s26r}) + r26r[39]);
		r27r[64:39]	<= r26r[64:39] ;
		r27r[4:0]	<= r26r[4:0] ;
		s27r <= s26r;

		// State: 28
		r28r[37:4]	<= ({r27r[38],r27r[36:4]}) + (({34{r27r[38]}}^{2'b00,s27r}) + r27r[38]);
		r28r[64:38]	<= r27r[64:38] ;
		r28r[3:0]	<= r27r[3:0] ;
		s28r <= s27r;

		// State: 29
		r29r[36:3]	<= ({r28r[37],r28r[35:3]}) + (({34{r28r[37]}}^{2'b00,s28r}) + r28r[37]);
		r29r[64:37]	<= r28r[64:37] ;
		r29r[2:0]	<= r28r[2:0] ;
		s29r <= s28r;

		// State: 30
		r30r[35:2]	<= ({r29r[36],r29r[34:2]}) + (({34{r29r[36]}}^{2'b00,s29r}) + r29r[36]);
		r30r[64:36]	<= r29r[64:36] ;
		r30r[1:0]	<= r29r[1:0] ;
		s30r <= s29r;

		// State: 31
		r31r[34:1]	<= ({r30r[35],r30r[33:1]}) + (({34{r30r[35]}}^{2'b00,s30r}) + r30r[35]);
		r31r[64:35]	<= r30r[64:35] ;
		r31r[0:0]	<= r30r[0:0] ;
		s31r <= s30r;

		// State: 32
		r32r[33:0]	<= ({r31r[34],r31r[32:0]}) + (({34{r31r[34]}}^{2'b00,s31r}) + r31r[34]);
		r32r[64:34]	<= r31r[64:34] ;

	end
end
assign DOUT = r32r[64:33];
endmodule
